// Author: Sriram Goparaju
// Date Created: 3/12/2022

module atpg (

	input 			clk,
	input 			rst,

	

);



endmodule // atpg